`ifndef M_get_radian
`define M_get_radian

module get_radian (
  input [4:0] address,
  output reg [21:0] data
);
    always @(*) begin
        case (address)
            5'd0:  data = 22'b1011010000000000000000;
            5'd1:  data = 22'b0110101001000010100111;
            5'd2:  data = 22'b0011100000100101000111;
            5'd3:  data = 22'b0001110010000000000001;
            5'd4:  data = 22'b0000111001001110001010;
            5'd5:  data = 22'b0000011100101000110111;
            5'd6:  data = 22'b0000001110010100101010;
            5'd7:  data = 22'b0000000111001010010110;
            5'd8:  data = 22'b0000000011100101001011;
            5'd9:  data = 22'b0000000001110010100101;
            5'd10: data = 22'b0000000000111001010010;
            5'd11: data = 22'b0000000000011100101001;
            5'd12: data = 22'b0000000000001110010100;
            5'd13: data = 22'b0000000000000111001010;
            5'd14: data = 22'b0000000000000011100101;
            5'd15: data = 22'b0000000000000001110010;
            5'd16: data = 22'b0000000000000000111001;
            5'd17: data = 22'b0000000000000000011100;
            5'd18: data = 22'b0000000000000000001110;
            5'd19: data = 22'b0000000000000000000111;
            5'd20: data = 22'b0000000000000000000011;
            5'd21: data = 22'b0000000000000000000001;
            default: data = 0;
        endcase
    end
endmodule

`endif